`timescale 1ns/1ps

`define max(a,b) {(a) > (b) ? (a) : (b)}
`define min(a,b) {(a) < (b) ? (a) : (b)}

/*WARNING: This memory assumes that the read port data width is bigger than the
write port data width and that they are multiples of eachother
*/
module iob_2p_assim_async_mem_r_big
	#( 
		parameter W_DATA_W = 16,
		parameter W_ADDR_W = 6,
		parameter R_DATA_W = 8,
		parameter R_ADDR_W = 7
	) 
	(
		//Inputs
	 input 			   wclk, //write clock
         input 			   w_en, //write enable
         input [W_DATA_W-1:0] 	   data_in, //Input data to write port
         input [W_ADDR_W-1:0] 	   w_addr, //address for write port
	 input 			   rclk, //read clock
         input [R_ADDR_W-1:0] 	   r_addr, //address for read port
         input 			   r_en,
        //Outputs
         output reg [R_DATA_W-1:0] data_out //output port
    );
	//local variables
	localparam maxADDR_W = `max(W_ADDR_W, R_ADDR_W);
	localparam maxDATA_W = `max(W_DATA_W, R_DATA_W);
	localparam minDATA_W = `min(W_DATA_W, R_DATA_W);
	localparam RATIO = maxDATA_W / minDATA_W;
	localparam log2RATIO = $clog2(RATIO);
	
	//memory declaration
	reg [minDATA_W-1:0] ram [2**maxADDR_W-1:0];
	
	integer i;
	reg [log2RATIO-1:0] lsbaddr;
	
	//writing to the RAM
	always@(posedge wclk)
		if (w_en)
			ram[gray2binW(w_addr, W_ADDR_W)] <= data_in;
	
	//reading from the RAM
	always@(posedge rclk) begin
		if (r_en) begin
			for (i = 0; i < RATIO; i = i+1) begin
				lsbaddr = i;
				data_out[(i+1)*minDATA_W-1 -: minDATA_W] <= ram[{gray2binR(r_addr, R_ADDR_W), lsbaddr}];
			end
		end
	end

      //convert gray to binary code - Write addresses
   function [W_ADDR_W-1:0] gray2binW;
      input reg [W_ADDR_W-1:0] gr;
      input integer 	       N;
      begin: g2b
	 reg [W_ADDR_W-1:0] bi;
	 integer 	    i;
	 
	 bi[N-1] = gr[N-1];
	 for (i=N-2;i>=0;i=i-1)
           bi[i] = gr[i] ^ bi[i+1];
	 
	 gray2binW = bi;
      end
   endfunction
   //convert gray to binary code - Read addresses
   function [R_ADDR_W-1:0] gray2binR;
      input reg [R_ADDR_W-1:0] gr;
      input integer 	       N;
      begin: g2b
	 reg [R_ADDR_W-1:0] bi;
	 integer 	    i;
	 
	 bi[N-1] = gr[N-1];
	 for (i=N-2;i>=0;i=i-1)
           bi[i] = gr[i] ^ bi[i+1];
	 
	 gray2binR = bi;
      end
   endfunction

endmodule   
