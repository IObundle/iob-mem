`define FIFO_DATA 0
`define FIFO_EMPTY 1
`define FIFO_FULL 2
`define FIFO_LEVEL_R 3
`define FIFO_LEVEL_W 4
`define FIFO_FLUSH 5
